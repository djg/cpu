//  ============================================================================
//  Copyright (C) 2018 Dan Glastonbury <dan.glastonbury@gmail.com>
//  ============================================================================

module cpu_counter(// ------ Inputs ------
                   clk_i,
                   rst_i,
                   // ------ Outputs -----
                   count_o
                   );

   //////////////////////////////////////////////////////
   // Inputs
   //////////////////////////////////////////////////////

   input clk_i;
   input rst_i;

   //////////////////////////////////////////////////////
   // Output
   //////////////////////////////////////////////////////

   output [3:0] count_o;

   //////////////////////////////////////////////////////
   // Interal nets and registers
   //////////////////////////////////////////////////////
   reg [3:0]    count_o;
   
   //////////////////////////////////////////////////////
   // Functions
   //////////////////////////////////////////////////////

   //////////////////////////////////////////////////////
   // Instantiations
   //////////////////////////////////////////////////////

   //////////////////////////////////////////////////////
   // Combinatorial Logic
   //////////////////////////////////////////////////////

   //////////////////////////////////////////////////////
   // Sequential Logic
   //////////////////////////////////////////////////////
   always @(posedge clk_i)
     begin
        if (rst_i == 1'b1) begin
           count_o <= 4'b0000;
        end
        else begin
           count_o <= count_o + 1;

        end
     end
   
   //////////////////////////////////////////////////////
   // Behavioural Logic
   //////////////////////////////////////////////////////
   
endmodule
